library ieee;
use ieee.std_logic_1164.all;

package myPackage is

	type ALU_operation is
		(ADDWF, ANDWF, COMF, DECF, INCF, SUBWF, ADDLW, ANDLW, SUBLW);

end myPackage;